module condlogic (
  clk,
  reset,
  Cond,
  ALUFlags,
  FlagW,
  PCS,
  RegW,
  MemW,
  PCSrc,
  RegWrite,
  MemWrite,
  Branch,
  BranchTakenE,
  BranchPredictor,
  FlagsE,
  FlagsNext
);
  input wire clk;
  input wire reset;
  input wire [3:0] Cond;
  input wire [3:0] ALUFlags;
  input wire [1:0] FlagW;
  input wire PCS;
  input wire RegW;
  input wire MemW;
  input wire Branch;
  input wire [3:0] FlagsE;
  output wire PCSrc;
  output wire RegWrite;
  output wire MemWrite;
  output wire BranchTakenE;
  output wire [3:0] FlagsNext;
  wire [1:0] FlagWrite;
  wire [3:0] Flags;
  wire CondEx;
  flopenr #(2) flagreg1 (
    .clk(clk),
    .reset(reset),
    .en(FlagWrite[1]),
    .d(ALUFlags[3:2]),
    .q(Flags[3:2])
  );
  flopenr #(2) flagreg0 (
    .clk(clk),
    .reset(reset),
    .en(FlagWrite[0]),
    .d(ALUFlags[1:0]),
    .q(Flags[1:0])
  );
  condcheck cc (
    .Cond(Cond),
    .Flags(Flags),
    .CondEx(CondEx)
  );
  assign FlagWrite = FlagW & {2{CondEx}};
  assign RegWrite = RegW & CondEx;
  assign MemWrite = MemW & CondEx;
  assign PCSrc = PCS & CondEx;
  assign BranchTakenE = Branch & CondEx;
  assign FlagsNext = Flags;

  output wire BranchPredictor;

  fsm BP1B (
    .clk(clk),
    .reset(reset),
    .ipt(BranchTakenE),
    .otpt(BranchPredictor)
  );
endmodule